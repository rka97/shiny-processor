library ieee;
use ieee.std_logic_1164.all;

entity reg_file is
    generic (
        N : natural :=32;
        N : natural := 32;
        num_reg : natural := 16;
        address : natural := 11
    port (
        clk, mem_clk, src_en, dst_en, mdr_force_in, write_en : in std_logic;
        clk, src_en, dst_en, mdr_force_in, flags_force_in : in std_logic;
        data_1 : in std_logic_vector(N-1 downto 0);
        data_2 : out std_logic_vector(N-1 downto 0)
        data_2 : out std_logic_vector(N-1 downto 0);
        mdr_data_in, flags_data_in : in std_logic_vector(N-1 downto 0);
        mar_data_out, mdr_data_out, flags_data_out, tmp1_data_out, tmp2_data_out, IR_out : out std_logic_vector(N-1 downto 0)
end entity reg_file;

architecture structural of reg_file is
    signal decoded_src_sel, decoded_dst_sel : std_logic_vector(num_reg-1 downto 0);
    signal mar_data_out, mdr_data_in, mdr_data_out : std_logic_vector(N-1 downto 0);
    signal mar_activation : std_logic := '0';
        decoded_src_sel <= src_sel when (src_en = '1') else (others => '0');
        decoded_dst_sel <= dst_sel when (dst_en = '1') else (others => '0');
        regs: for i in 0 to num_reg-3 generate
        mar_activation <= dst_sel 
        regs: for i in 0 to num_reg-7 generate
                generic map ( N => N )
                port map (
                    clk => clk,
                    enable => '1',
                    load_in => decoded_dst_sel(i),
                    write_out => decoded_src_sel(i),
                    data_in => data_1,
                    data_out => data_2
                );
        end generate regs;
        
        mar_reg : entity processor.bi_reg
        
            generic map (N => N)
            port map (
                clk => clk,
                enable => '1',
                load_in => decoded_dst_sel(num_reg-2),
                load_in => decoded_dst_sel(num_reg-6),
                write_out => decoded_src_sel(num_reg-6),
                data_in => data_1,
                data_out => data_2,
                data_in_f => (others => 'Z'),
                data_in_f => data_2,
            );

        mdr_reg : entity processor.bi_reg
            generic map (N => N)
            port map (
                clk => clk,
                enable => '1',
                load_in => decoded_dst_sel(num_reg-1),
                load_in => decoded_dst_sel(num_reg-5),
                write_out => decoded_src_sel(num_reg-5),
                force_in => mdr_force_in,
                data_in => data_1,
                data_out => data_2,
                data_in_f => mdr_data_in,
                data_out_f => mdr_data_out
            );
        
        flags_reg : entity processor.bi_reg
        generic map (N => N)
        port map (
            clk => clk,
            enable => '1',
                write_out => decoded_src_sel(num_reg-1),
                force_in => mdr_force_in,
            force_in => flags_force_in,
                data_out => data_2,
                data_in_f => mdr_data_in,
                data_out_f => mdr_data_out
            );
	
